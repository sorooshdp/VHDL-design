
entity four_to_sixteen is
end four_to_sixteen;

--}} End of automatically maintained section

architecture four_to_sixteen of four_to_sixteen is
begin

	 -- enter your statements here --

end four_to_sixteen;
